module not_func (
    input [7:0] in1,
    input [7:0] in2,
    output [7:0] out
);
    // Implement not!
    assign out = ~in1;
endmodule

module or_tb(
)
endmodule